`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// ECE369 - Computer Architecture
// 
// Module - SignExtension.v
// Description - Sign extension module.
////////////////////////////////////////////////////////////////////////////////
module SignExtension(in, ZeroExtend, out);

    /* A 16-Bit input word */
    input [15:0] in;
    
    /* A 32-Bit output word */
    output reg [31:0] out;
    
    /* Fill in the implementation here ... */
    input ZeroExtend;
    always @(*) begin
        if(ZeroExtend) begin
            out = {16'h0000, in};
        end
        else begin
            if(in[15] == 1) begin
                out = {16'hFFFF, in};
            end
            else begin
                out = {16'h0000, in};
            end
        end
    end
endmodule
