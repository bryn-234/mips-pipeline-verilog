`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory 1
// Module - ProgramCounter_tb.v
// Description - Test the 'ProgramCounter.v' module.
////////////////////////////////////////////////////////////////////////////////

module ProgramCounter_tb(); 

	reg [31:0] Address;
	reg Reset, Clk;

	wire [31:0] PCResult;

    ProgramCounter u0(
        .Address(Address), 
        .PCResult(PCResult), 
        .Reset(Reset), 
        .Clk(Clk)
    );

	initial begin
		Clk <= 1'b0;
		forever #10 Clk <= ~Clk;
	end

	initial begin
	
    /* Please fill in the implementation here... */
	   @(posedge Clk)
	   Address <= 32'd0;
	   #10
	   
	   @(posedge Clk)
	   Address <= 32'd4;
	   #10
	   
	   @(posedge Clk)
	   Address <= 32'd8;
	   #10
	   
	   @(posedge Clk)
	   Address <= 32'd12;
	   #10
	   
	   @(posedge Clk)
	   Address <= 32'd16;
	   #10
	   
	   @(posedge Clk)
	   Address <= 32'd20;
	   
	end

endmodule

